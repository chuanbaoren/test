module fifo()
