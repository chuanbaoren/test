module fifo()
222222
